//-----------------------------------------------------
// File Name   : alucodes.sv
// Function    : pMIPS ALU function code definiRons
// Author:  rz
// Last rev. 24/04/2024
//-----------------------------------------------------

//`define RNOP    3'b000
`define RADD    1'b0

`define RMUL    1'b1